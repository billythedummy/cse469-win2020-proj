/*
module mux
    #(parameter inputs=4,
        parameter width=8)
    (out, ); 

endmodule
*/  