module idec () //instruction decoder

endmodule