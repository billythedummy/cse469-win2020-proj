module regfile ();
    
endmodule